`timescale 1ns / 1ps
module boolean_expression(input a, b, c, output y);
assign y = (a & b) | (~a & c);
endmodule


module boolean_expression(

    );
endmodule
