`timescale 1ns / 1ps
module boolean_expression_tb;
reg a, b, c;
wire y;

boolean_expression uut(a, b, c, y);

initial begin
$monitor("Time=%0t | a=%b b=%b c=%b | y=%b", $time, a, b, c, y);
a=0; b=0; c=0;
#10 a=0; b=0; c=1;
#10 a=0; b=1; c=0;
#10 a=0; b=1; c=1;
#10 a=1; b=0; c=0;
#10 a=1; b=0; c=1;
#10 a=1; b=1; c=0;
#10 a=1; b=1; c=1;
#10 $finish;
end
endmodule

//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.11.2025 21:19:36
// Design Name: 
// Module Name: boolean_expression_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module boolean_expression_tb(

    );
endmodule
